--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use WORK.st7735r_p_package.ALL;

package st7735r_p_store_image_data is

	constant R_EDGE : std_logic := '1';
	constant F_EDGE : std_logic := '0';
	subtype byte is std_logic_vector(0 to BYTE_SIZE-1);
	constant Xs : std_logic_vector(0 to BYTE_SIZE - 1) := (others => 'U');
	
	type states1 is (idle,start_cs,ck_event,ck_event_increment,stop_cs);
	shared variable state1 : states1;
	type states2 is (idle,pattern1,pattern2,pattern3,start,stop);
	shared variable state2 : states2;

	shared variable data_temp_index : integer;

	shared variable do_temp : byte;

	shared variable done : std_logic;
	shared variable do_data : byte;

	function vec2str(vec: std_logic_vector) return string;

	procedure spi_get_byte (
		signal i_clock : in std_logic;
		signal i_reset : in std_logic;
		signal cs : in std_logic;
		signal do : in std_logic;
		signal ck : in std_logic;
		variable done : out std_logic;
		variable do_data : inout byte
	);

	procedure st7735r_store_image_fsm (
		signal i_clock : in std_logic;
		signal i_reset : in std_logic;
		signal cs : in std_logic;
		signal do : in std_logic;
		signal ck : in std_logic
	);

end st7735r_p_store_image_data;

package body st7735r_p_store_image_data is

	procedure spi_get_byte (
		signal i_clock : in std_logic;
		signal i_reset : in std_logic;
		signal cs : in std_logic;
		signal do : in std_logic;
		signal ck : in std_logic;
		variable done : out std_logic;
		variable do_data : inout byte -- XXX default out, inout for report
	) is
	begin
		if (i_reset = '1') then
			state1 := idle;
			data_temp_index := 0;
			do_temp := (others => '0');
			done := '0';
		elsif (rising_edge(i_clock)) then
			case (state1) is
				when idle =>
					state1 := start_cs;
					data_temp_index := 0;
					do_temp := (others => '0');
					done := '0';
				when start_cs =>
					if (cs = '0') then
						state1 := ck_event;
--						report "spi_get_byte cs = '0'" severity note;
					else
						state1 := start_cs;
					end if;
				when ck_event =>
					if (ck = R_EDGE) then
						state1 := ck_event_increment;
						do_temp(data_temp_index) := do;
					else
						state1 := ck_event;
					end if;
				when ck_event_increment =>
					if (data_temp_index = BYTE_SIZE - 1) then
						state1 := stop_cs;
					else
						state1 := ck_event;
						data_temp_index := data_temp_index + 1;
					end if;
				when stop_cs =>
					if (cs = '1') then
						state1 := idle;
						do_data := do_temp;
						done := '1';
--						report "spi_get_byte cs = '1'" severity note;
						report "spi_get_byte do_data = " & vec2str(do_data) severity note;
					elsif (cs = '0') then
						state1 := stop_cs;
					end if;
			end case;
		end if;
	end procedure spi_get_byte;

	procedure st7735r_store_image_fsm (
		signal i_clock : in std_logic;
		signal i_reset : in std_logic;
		signal cs : in std_logic;
		signal do : in std_logic;
		signal ck : in std_logic
	) is
--		variable do_data : byte;
--		variable state : states; -- XXX must stay variable, "Signal declaration is not allowed in a subprogram"
--		variable done : std_logic;
	begin
		if (i_reset = '1') then
			state2 := idle;
--			do_data <= (others => 'U');
--			spi_get_byte(i_clock,i_reset,cs,do,ck,do_data,done);
		elsif (rising_edge(i_clock)) then
			case (state2) is
				when idle =>
					if (cs = '1') then
						state2 := idle;
					else
						state2 := pattern1;
					end if;
				when pattern1 =>
					if (do_data = x"2b") then
						state2 := pattern2;
					else
						state2 := pattern1;
					end if;
				when pattern2 =>
					if (do_data = x"2a") then
						state2 := pattern3;
					else
						state2 := pattern2;
					end if;
				when pattern3 =>
					if (do_data = x"2c") then
						state2 := start;
					else
						state2 := pattern3;
					end if;
				when start =>
					state2 := stop;
					report "asd" severity note;
				when stop =>
					state2 := idle;
			end case;
		end if;
					spi_get_byte(i_clock,i_reset,cs,do,ck,done,do_data);

	end procedure st7735r_store_image_fsm;

	function vec2str(vec: std_logic_vector) return string is
		variable result: string(0 to vec'right);
	begin
		for i in vec'range loop
			if (vec(i) = '1') then
				result(i) := '1';
			elsif (vec(i) = '0') then
				result(i) := '0';
			elsif (vec(i) = 'X') then
				result(i) := 'X';
			elsif (vec(i) = 'U') then
				result(i) := 'U';
			else
				result(i) := '?';
			end if;
		end loop;
		return result;
	end;

--			assert (data_rom(data_rom_index) = data_temp) report "FAIL : (" & integer'image(data_rom_index) & ") " & vec2str(data_temp) & " expect " & vec2str(data_rom(data_rom_index)) severity note;
--			assert (data_rom(data_rom_index) /= data_temp) report "OK   : (" & integer'image(data_rom_index) & ") " & vec2str(data_temp) & " equals " & vec2str(data_rom(data_rom_index)) severity note;
--			data_temp_index := 0;
--			if (data_rom_index = data_size - 1) then
--				data_rom_index := 0;
--				assert (false) report "=== END TEST ===" severity note;
--			else
--				if (data_temp /= Xs) then -- XXX omit first undefined/uninitialized
--					data_rom_index := data_rom_index + 1;
--				end if;
--			end if;

end st7735r_p_store_image_data;
