entity n2_core_pll_pad_cluster_cust is
port(
vdd_hv15 : in bit;
pll_sys_clk : in bit_vector(1 downto 0)
);
end entity n2_core_pll_pad_cluster_cust;
architecture arch of n2_core_pll_pad_cluster_cust is
--supply1 vdd ;
begin
end architecture arch; 

