----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:07:54 10/27/2020 
-- Design Name: 
-- Module Name:    memory1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity memory1 is
Generic (
WIDTH : integer := 128;
HEIGHT : integer := 32;
W_BITS : integer := 7;
H_BITS : integer := 5);
Port (
i_clk : in std_logic;
i_x : in std_logic_vector(W_BITS-1 downto 0);
i_y : in std_logic_vector(H_BITS-1 downto 0);
o_bit : out std_logic_vector(0 downto 0));
end memory1;

architecture Behavioral of memory1 is
	type array1 is array(0 to WIDTH-1) of std_logic_vector(0 to HEIGHT-1);
	
-- https://www.conwaylife.com/patterns/gosperglidergun.cells
-- !Name: Gosper glider gun
-- !Author: Bill Gosper
-- !The first known gun and the first known finite pattern with unbounded growth.
-- !www.conwaylife.com/wiki/index.php?title=Gosper_glider_gun
-- ........................O
-- ......................O.O
-- ............OO......OO............OO
-- ...........O...O....OO............OO
-- OO........O.....O...OO
-- OO........O...O.OO....O.O
-- ..........O.....O.......O
-- ...........O...O
-- ............OO

	signal m1 : array1 :=
	(
		("00000000000000000000000010000000"),
		("00000000000000000000001010000000"),
		("00000000000011000000110000000000"),
		("00000000000100010000110000000000"),
		("11000000001000001000110000000000"),
		("11000000001000101100001010000000"),
		("00000000001000001000000010000000"),
		("00000000000100010000000000000000"),
		("00000000000011000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000"),
		("00000000000000000000000000000000")
	);
begin
	o_bit(0) <= m1(to_integer(unsigned(i_x)))(to_integer(unsigned(i_y)));
end Behavioral;
