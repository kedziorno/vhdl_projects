--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   11:39:28 04/19/2021
-- Design Name:   
-- Module Name:   /home/user/workspace/vhdl_projects/vhdl_primitive/tb_pwm_generator.vhd
-- Project Name:  vhdl_primitive
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: PWM_generator
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
USE ieee.numeric_std.ALL;

ENTITY tb_pwm_generator IS
END tb_pwm_generator;

ARCHITECTURE behavior OF tb_pwm_generator IS

constant N : integer := 4;

-- Component Declaration for the Unit Under Test (UUT)
COMPONENT PWM_generator
GENERIC(N : integer);
PORT(
i_clock : IN  std_logic;
i_reset : IN  std_logic;
i_data : IN  std_logic_vector(N-1 downto 0);
o_pwm : OUT  std_logic
);
END COMPONENT;

--Inputs
signal i_clock : std_logic := '0';
signal i_reset : std_logic := '0';
signal i_data : std_logic_vector(N-1 downto 0) := (others => '0');

--Outputs
signal o_pwm : std_logic;

-- Clock period definitions
constant i_clock_period : time := 20 ns;

BEGIN

-- Instantiate the Unit Under Test (UUT)
uut: PWM_generator 
GENERIC MAP (N => N)
PORT MAP (
i_clock => i_clock,
i_reset => i_reset,
i_data => i_data,
o_pwm => o_pwm
);

-- Clock process definitions
i_clock_process :process
begin
i_clock <= '0';
wait for i_clock_period/2;
i_clock <= '1';
wait for i_clock_period/2;
end process;

-- Stimulus process
stim_proc: process
begin
-- hold reset state for 100 ns.
i_reset <= '1';
wait for 100 ns;
i_reset <= '0';
wait for i_clock_period*10;
-- insert stimulus here
l0 : for i in 0 to (2**N)-1 loop
i_data <= std_logic_vector(to_unsigned(i,N));
wait for i_clock_period*(2**N)*2;
end loop l0;
i_data <= std_logic_vector(to_unsigned(0,N));
wait for i_clock_period*(2**N)*2;
wait;
end process;

END;
