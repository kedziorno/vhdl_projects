----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:47:31 08/21/2020 
-- Design Name: 
-- Module Name:    power_on - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use WORK.p_constants1.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
use ieee.std_logic_unsigned.all;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity power_on is 
port (
	i_clock : in std_logic;
	i_reset : in std_logic;
	o_sda : out std_logic;
	o_scl : out std_logic
);
end power_on;

architecture Behavioral of power_on is

	COMPONENT my_i2c IS
	GENERIC (
		BOARD_CLOCK : INTEGER := G_BOARD_CLOCK;
		BUS_CLOCK : INTEGER := G_BUS_CLOCK;
		SEQUENCE_LENGTH : INTEGER := 1
	);
	PORT (
		i_clock : in std_logic;
		i_reset : in std_logic;
		i_slave_address : std_logic_vector(G_SLAVE_ADDRESS_SIZE-1 downto 0);
		i_bytes_to_send : array_byte_sequence(0 to SEQUENCE_LENGTH-1);
		i_enable : in std_logic;
		o_busy : out std_logic;
		o_sda : out std_logic;
		o_scl : out std_logic
	);
	END COMPONENT my_i2c;

begin

	my_i2c_entity : my_i2c
	GENERIC MAP (
		BOARD_CLOCK => G_BOARD_CLOCK,
		BUS_CLOCK => G_BUS_CLOCK,
		SEQUENCE_LENGTH => BYTES_SEQUENCE_LENGTH
	)
	PORT MAP (
		i_clock => i_clock,
		i_reset => i_reset,
		i_slave_address => "0111100",
		i_bytes_to_send => sequence,
		i_enable => '1',
		o_busy => open,
		o_sda => o_sda,
		o_scl => o_scl
	);

end Behavioral;
