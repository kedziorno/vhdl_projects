library IEEE;
use IEEE.STD_LOGIC_1164.all;

package p_globals is
end p_globals;

package body p_globals is
end p_globals;

