----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:11:00 11/28/2020
-- Design Name: 
-- Module Name:    /home/user/workspace/vhdl_projects/memorymodule/memorymodule.vhd
-- Project Name:   memorymodule
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use WORK.p_memory_content.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity memorymodule_bram is
Port (
i_clock : in std_logic;
i_enable : in std_logic;
i_write : in std_logic;
i_read : in std_logic;
o_busy : out std_logic;
i_MemAdr : in MemoryAddress;
i_MemDB : in MemoryDataByte;
o_MemDB : out MemoryDataByte;
o_MemOE : out std_logic;
o_MemWR : out std_logic;
o_RamAdv : out std_logic;
o_RamCS : out std_logic;
o_RamCRE : out std_logic;
o_RamLB : out std_logic;
o_RamUB : out std_logic;
i_RamWait : in std_logic;
o_RamClk : out std_logic;
o_MemAdr : out MemoryAddress;
io_MemDB : inout MemoryDataByte
);
end memorymodule_bram;

architecture Behavioral of memorymodule_bram is

type state is (
idle,
start,
write_setup,
read_setup,
write_enable,
wait1,
write_disable,
stop,
read1,
wait2
);
signal cstate : state;

signal MemOE : std_logic;
signal MemWR : std_logic;
signal RamAdv : std_logic;
signal RamCS : std_logic;
signal RamLB : std_logic;
signal RamCRE : std_logic;
signal RamUB : std_logic;
signal RamClk : std_logic;
signal MemAdr : MemoryAddress;
signal MemDB : MemoryDataByte;

signal RAMB36_S18_DO,RAMB36_S18_DI : std_logic_vector(15 downto 0);
signal RAMB36_S18_DOP,RAMB36_S18_DIP : std_logic_vector(1 downto 0);
signal RAMB36_S18_ADDR : std_logic_vector(9 downto 0);
signal RAMB36_S18_CLK,RAMB36_S18_EN,RAMB36_S18_SSR,RAMB36_S18_WE : std_logic;

begin

--MemAdr <= i_MemAdr when (RamCS = '0' and (MemWR = '0' or MemOE = '0')) else (others => 'Z');
--o_MemDB <= io_MemDB when (cstate = idle) else (others => 'Z');
--io_MemDB <= i_MemDB when (RamCS = '0' and MemWR = '0') else (others => 'Z');

RAMB36_S18_ADDR(9 downto 0) <= i_MemAdr(10 downto 1) when (RamCS = '0' and (MemWR = '0' or MemOE = '0')) else (others => 'Z');
io_MemDB <= RAMB36_S18_DO when (cstate = idle) else (others => 'Z');
--io_MemDB <= RAMB36_S18_DO when (cstate = idle or cstate = start or cstate = read_setup or cstate = read1 or cstate = wait2) else (others => 'Z');
o_MemDB <= RAMB36_S18_DO when (RamCS = '0' and MemOE = '0') else (others => 'Z');
RAMB36_S18_DI <= i_MemDB when (RamCS = '0' and MemWR = '0') else (others => 'Z');
RAMB36_S18_CLK <= i_clock;
RAMB36_S18_EN <= not RamCS;
--RAMB36_S18_EN <= '1';
RAMB36_S18_WE <= not MemWR;
RAMB36_S18_SSR <= '0';

o_MemAdr <= MemAdr;
o_RamCS <= RamCS;
o_MemOE <= MemOE;
o_MemWR <= MemWR;

o_RamAdv <= RamAdv;
o_RamClk <= RamClk;
o_RamCRE <= RamCRE;
o_RamLB <= RamLB;
o_RamUB <= RamUB;

RamAdv <= '0';
RamClk <= '0';
RamCRE <= '0';
RamLB <= '0';
RamUB <= '0';

p0 : process (i_clock) is
	constant cw : integer := 6;
	variable w : integer range 0 to cw := 0;
	variable t : std_logic_vector(G_MemoryData-1 downto 0);
	variable tz : std_logic_vector(G_MemoryData-1 downto 0) := (others => 'Z');
begin
	if (rising_edge(i_clock)) then
		if (w > 0) then
			w := w - 1;
		end if;
		case cstate is
			when idle =>
				if (i_enable = '1') then
					cstate <= start; -- XXX check CSb
				else
					cstate <= idle;
				end if;
			when start =>
				if (i_write = '1') then
					cstate <= write_setup;
				elsif (i_read = '1') then
					cstate <= read_setup;
				else
					cstate <= start;
				end if;
				RamCS <= '1';
				MemWR <= '1';
				MemOE <= '1';
			when write_setup =>
				if (w = 0) then
					cstate <= write_enable;
					o_busy <= '1';
					MemOE <= '1';
				else
					cstate <= write_setup;
				end if;
			when write_enable =>
				cstate <= wait1;
				MemWR <= '0';
				RamCS <= '0';
				w := cw;
			when wait1 =>
				if (w = 0) then
					cstate <= write_disable;
				else
					cstate <= wait1;
				end if;
			when write_disable =>
				cstate <= stop;
				RamCS <= '1';
				MemWR <= '1';
			when read_setup =>
				if (w = 0) then
					cstate <= read1;
					RamCS <= '0';
					MemOE <= '0';
					o_busy <= '1';
				else
					cstate <= read_setup;
				end if;
			when read1 =>
				cstate <= wait2;
				w := cw;
			when wait2 =>
				if (w = 0) then
					cstate <= stop;
				else
					cstate <= wait2;
				end if;
			when stop =>
				cstate <= idle;
				o_busy <= '0';
				RamCS <= '1';
				MemOE <= '1';
			when others => null;
		end case;
	end if;
end process p0;

-- RAMB16_S18: 1k x 16 + 2 Parity bits Single-Port RAM
-- Spartan-3E
-- Xilinx HDL Libraries Guide, version 14.5
RAMB16_S18_inst : RAMB16_S18
generic map (
INIT => X"00000", -- Value of output RAM registers at startup
SRVAL => X"00000", -- Output value upon SSR assertion
WRITE_MODE => "NO_CHANGE", -- WRITE_FIRST, READ_FIRST or NO_CHANGE
-- The following INIT_xx declarations specify the intial contents of the RAM
-- Address 0 to 255
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- Address 256 to 511
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- Address 512 to 767
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- Address 768 to 1023
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- The next set of INITP_xx are for the parity bits
-- Address 0 to 255
INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- Address 256 to 511
INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- Address 512 to 767
INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- Address 768 to 1023
INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
port map (
DO => RAMB36_S18_DO, -- 16-bit Data Output
DOP => RAMB36_S18_DOP, -- 2-bit parity Output
ADDR => RAMB36_S18_ADDR, -- 10-bit Address Input
CLK => RAMB36_S18_CLK, -- Clock
DI => RAMB36_S18_DI, -- 16-bit Data Input
DIP => RAMB36_S18_DIP, -- 2-bit parity Input
EN => RAMB36_S18_EN, -- RAM Enable Input
SSR => RAMB36_S18_SSR, -- Synchronous Set/Reset Input
WE => RAMB36_S18_WE -- Write Enable Input
);

end Behavioral;
