library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity glcdfont is
port (
signal i_clk : in std_logic;
signal i_reset : in std_logic;
signal i_index : in std_logic_vector(10 downto 0);
signal o_character : out std_logic_vector(7 downto 0)
);
end entity glcdfont;

architecture behavioral_glcdfont of glcdfont is

constant NUMBER_GLCDFONTC : natural := 1275;
type ARRAY_GLCDFONTC is array (0 to NUMBER_GLCDFONTC-1) of std_logic_vector(7 downto 0);
constant GLCDFONTC : ARRAY_GLCDFONTC :=
(

	 -- 0:    0x00, 0x00, 0x00, 0x00, 0x00,   
	x"00",
	x"00",
	x"00",
	x"00",
	x"00",

	 -- 5:	0x3E, 0x5B, 0x4F, 0x5B, 0x3E, 	
	x"3E",
	x"5B",
	x"4F",
	x"5B",
	x"3E",

	 -- 10:	0x3E, 0x6B, 0x4F, 0x6B, 0x3E, 	
	x"3E",
	x"6B",
	x"4F",
	x"6B",
	x"3E",

	 -- 15:	0x1C, 0x3E, 0x7C, 0x3E, 0x1C, 
	x"1C",
	x"3E",
	x"7C",
	x"3E",
	x"1C",

	 -- 20:	0x18, 0x3C, 0x7E, 0x3C, 0x18, 
	x"18",
	x"3C",
	x"7E",
	x"3C",
	x"18",

	 -- 25:	0x1C, 0x57, 0x7D, 0x57, 0x1C, 
	x"1C",
	x"57",
	x"7D",
	x"57",
	x"1C",

	 -- 30:	0x1C, 0x5E, 0x7F, 0x5E, 0x1C, 
	x"1C",
	x"5E",
	x"7F",
	x"5E",
	x"1C",

	 -- 35:	0x00, 0x18, 0x3C, 0x18, 0x00, 
	x"00",
	x"18",
	x"3C",
	x"18",
	x"00",

	 -- 40:	0xFF, 0xE7, 0xC3, 0xE7, 0xFF, 
	x"FF",
	x"E7",
	x"C3",
	x"E7",
	x"FF",

	 -- 45:	0x00, 0x18, 0x24, 0x18, 0x00, 
	x"00",
	x"18",
	x"24",
	x"18",
	x"00",

	 -- 50:	0xFF, 0xE7, 0xDB, 0xE7, 0xFF, 
	x"FF",
	x"E7",
	x"DB",
	x"E7",
	x"FF",

	 -- 55:	0x30, 0x48, 0x3A, 0x06, 0x0E, 
	x"30",
	x"48",
	x"3A",
	x"06",
	x"0E",

	 -- 60:	0x26, 0x29, 0x79, 0x29, 0x26, 
	x"26",
	x"29",
	x"79",
	x"29",
	x"26",

	 -- 65:	0x40, 0x7F, 0x05, 0x05, 0x07, 
	x"40",
	x"7F",
	x"05",
	x"05",
	x"07",

	 -- 70:	0x40, 0x7F, 0x05, 0x25, 0x3F, 
	x"40",
	x"7F",
	x"05",
	x"25",
	x"3F",

	 -- 75:	0x5A, 0x3C, 0xE7, 0x3C, 0x5A, 
	x"5A",
	x"3C",
	x"E7",
	x"3C",
	x"5A",

	 -- 80:	0x7F, 0x3E, 0x1C, 0x1C, 0x08, 
	x"7F",
	x"3E",
	x"1C",
	x"1C",
	x"08",

	 -- 85:	0x08, 0x1C, 0x1C, 0x3E, 0x7F, 
	x"08",
	x"1C",
	x"1C",
	x"3E",
	x"7F",

	 -- 90:	0x14, 0x22, 0x7F, 0x22, 0x14, 
	x"14",
	x"22",
	x"7F",
	x"22",
	x"14",

	 -- 95:	0x5F, 0x5F, 0x00, 0x5F, 0x5F, 
	x"5F",
	x"5F",
	x"00",
	x"5F",
	x"5F",

	 -- 100:	0x06, 0x09, 0x7F, 0x01, 0x7F, 
	x"06",
	x"09",
	x"7F",
	x"01",
	x"7F",

	 -- 105:	0x00, 0x66, 0x89, 0x95, 0x6A, 
	x"00",
	x"66",
	x"89",
	x"95",
	x"6A",

	 -- 110:	0x60, 0x60, 0x60, 0x60, 0x60, 
	x"60",
	x"60",
	x"60",
	x"60",
	x"60",

	 -- 115:	0x94, 0xA2, 0xFF, 0xA2, 0x94, 
	x"94",
	x"A2",
	x"FF",
	x"A2",
	x"94",

	 -- 120:	0x08, 0x04, 0x7E, 0x04, 0x08, 
	x"08",
	x"04",
	x"7E",
	x"04",
	x"08",

	 -- 125:	0x10, 0x20, 0x7E, 0x20, 0x10, 
	x"10",
	x"20",
	x"7E",
	x"20",
	x"10",

	 -- 130:	0x08, 0x08, 0x2A, 0x1C, 0x08, 
	x"08",
	x"08",
	x"2A",
	x"1C",
	x"08",

	 -- 135:	0x08, 0x1C, 0x2A, 0x08, 0x08, 
	x"08",
	x"1C",
	x"2A",
	x"08",
	x"08",

	 -- 140:	0x1E, 0x10, 0x10, 0x10, 0x10, 
	x"1E",
	x"10",
	x"10",
	x"10",
	x"10",

	 -- 145:	0x0C, 0x1E, 0x0C, 0x1E, 0x0C, 
	x"0C",
	x"1E",
	x"0C",
	x"1E",
	x"0C",

	 -- 150:	0x30, 0x38, 0x3E, 0x38, 0x30, 
	x"30",
	x"38",
	x"3E",
	x"38",
	x"30",

	 -- 155:	0x06, 0x0E, 0x3E, 0x0E, 0x06, 
	x"06",
	x"0E",
	x"3E",
	x"0E",
	x"06",

	 -- 160:	0x00, 0x00, 0x00, 0x00, 0x00, 
	x"00",
	x"00",
	x"00",
	x"00",
	x"00",

	 -- 165:	0x00, 0x00, 0x5F, 0x00, 0x00, 
	x"00",
	x"00",
	x"5F",
	x"00",
	x"00",

	 -- 170:	0x00, 0x07, 0x00, 0x07, 0x00, 
	x"00",
	x"07",
	x"00",
	x"07",
	x"00",

	 -- 175:	0x14, 0x7F, 0x14, 0x7F, 0x14, 
	x"14",
	x"7F",
	x"14",
	x"7F",
	x"14",

	 -- 180:	0x24, 0x2A, 0x7F, 0x2A, 0x12, 
	x"24",
	x"2A",
	x"7F",
	x"2A",
	x"12",

	 -- 185:	0x23, 0x13, 0x08, 0x64, 0x62, 
	x"23",
	x"13",
	x"08",
	x"64",
	x"62",

	 -- 190:	0x36, 0x49, 0x56, 0x20, 0x50, 
	x"36",
	x"49",
	x"56",
	x"20",
	x"50",

	 -- 195:	0x00, 0x08, 0x07, 0x03, 0x00, 
	x"00",
	x"08",
	x"07",
	x"03",
	x"00",

	 -- 200:	0x00, 0x1C, 0x22, 0x41, 0x00, 
	x"00",
	x"1C",
	x"22",
	x"41",
	x"00",

	 -- 205:	0x00, 0x41, 0x22, 0x1C, 0x00, 
	x"00",
	x"41",
	x"22",
	x"1C",
	x"00",

	 -- 210:	0x2A, 0x1C, 0x7F, 0x1C, 0x2A, 
	x"2A",
	x"1C",
	x"7F",
	x"1C",
	x"2A",

	 -- 215:	0x08, 0x08, 0x3E, 0x08, 0x08, 
	x"08",
	x"08",
	x"3E",
	x"08",
	x"08",

	 -- 220:	0x00, 0x80, 0x70, 0x30, 0x00, 
	x"00",
	x"80",
	x"70",
	x"30",
	x"00",

	 -- 225:	0x08, 0x08, 0x08, 0x08, 0x08, 
	x"08",
	x"08",
	x"08",
	x"08",
	x"08",

	 -- 230:	0x00, 0x00, 0x60, 0x60, 0x00, 
	x"00",
	x"00",
	x"60",
	x"60",
	x"00",

	 -- 235:	0x20, 0x10, 0x08, 0x04, 0x02, 
	x"20",
	x"10",
	x"08",
	x"04",
	x"02",

	 -- 240:	0x3E, 0x51, 0x49, 0x45, 0x3E, 
	x"3E",
	x"51",
	x"49",
	x"45",
	x"3E",

	 -- 245:	0x00, 0x42, 0x7F, 0x40, 0x00, 
	x"00",
	x"42",
	x"7F",
	x"40",
	x"00",

	 -- 250:	0x72, 0x49, 0x49, 0x49, 0x46, 
	x"72",
	x"49",
	x"49",
	x"49",
	x"46",

	 -- 255:	0x21, 0x41, 0x49, 0x4D, 0x33, 
	x"21",
	x"41",
	x"49",
	x"4D",
	x"33",

	 -- 260:	0x18, 0x14, 0x12, 0x7F, 0x10, 
	x"18",
	x"14",
	x"12",
	x"7F",
	x"10",

	 -- 265:	0x27, 0x45, 0x45, 0x45, 0x39, 
	x"27",
	x"45",
	x"45",
	x"45",
	x"39",

	 -- 270:	0x3C, 0x4A, 0x49, 0x49, 0x31, 
	x"3C",
	x"4A",
	x"49",
	x"49",
	x"31",

	 -- 275:	0x41, 0x21, 0x11, 0x09, 0x07, 
	x"41",
	x"21",
	x"11",
	x"09",
	x"07",

	 -- 280:	0x36, 0x49, 0x49, 0x49, 0x36, 
	x"36",
	x"49",
	x"49",
	x"49",
	x"36",

	 -- 285:	0x46, 0x49, 0x49, 0x29, 0x1E, 
	x"46",
	x"49",
	x"49",
	x"29",
	x"1E",

	 -- 290:	0x00, 0x00, 0x14, 0x00, 0x00, 
	x"00",
	x"00",
	x"14",
	x"00",
	x"00",

	 -- 295:	0x00, 0x40, 0x34, 0x00, 0x00, 
	x"00",
	x"40",
	x"34",
	x"00",
	x"00",

	 -- 300:	0x00, 0x08, 0x14, 0x22, 0x41, 
	x"00",
	x"08",
	x"14",
	x"22",
	x"41",

	 -- 305:	0x14, 0x14, 0x14, 0x14, 0x14, 
	x"14",
	x"14",
	x"14",
	x"14",
	x"14",

	 -- 310:	0x00, 0x41, 0x22, 0x14, 0x08, 
	x"00",
	x"41",
	x"22",
	x"14",
	x"08",

	 -- 315:	0x02, 0x01, 0x59, 0x09, 0x06, 
	x"02",
	x"01",
	x"59",
	x"09",
	x"06",

	 -- 320:	0x3E, 0x41, 0x5D, 0x59, 0x4E, 
	x"3E",
	x"41",
	x"5D",
	x"59",
	x"4E",

	 -- 325:	0x7C, 0x12, 0x11, 0x12, 0x7C, 
	x"7C",
	x"12",
	x"11",
	x"12",
	x"7C",

	 -- 330:	0x7F, 0x49, 0x49, 0x49, 0x36, 
	x"7F",
	x"49",
	x"49",
	x"49",
	x"36",

	 -- 335:	0x3E, 0x41, 0x41, 0x41, 0x22, 
	x"3E",
	x"41",
	x"41",
	x"41",
	x"22",

	 -- 340:	0x7F, 0x41, 0x41, 0x41, 0x3E, 
	x"7F",
	x"41",
	x"41",
	x"41",
	x"3E",

	 -- 345:	0x7F, 0x49, 0x49, 0x49, 0x41, 
	x"7F",
	x"49",
	x"49",
	x"49",
	x"41",

	 -- 350:	0x7F, 0x09, 0x09, 0x09, 0x01, 
	x"7F",
	x"09",
	x"09",
	x"09",
	x"01",

	 -- 355:	0x3E, 0x41, 0x41, 0x51, 0x73, 
	x"3E",
	x"41",
	x"41",
	x"51",
	x"73",

	 -- 360:	0x7F, 0x08, 0x08, 0x08, 0x7F, 
	x"7F",
	x"08",
	x"08",
	x"08",
	x"7F",

	 -- 365:	0x00, 0x41, 0x7F, 0x41, 0x00, 
	x"00",
	x"41",
	x"7F",
	x"41",
	x"00",

	 -- 370:	0x20, 0x40, 0x41, 0x3F, 0x01, 
	x"20",
	x"40",
	x"41",
	x"3F",
	x"01",

	 -- 375:	0x7F, 0x08, 0x14, 0x22, 0x41, 
	x"7F",
	x"08",
	x"14",
	x"22",
	x"41",

	 -- 380:	0x7F, 0x40, 0x40, 0x40, 0x40, 
	x"7F",
	x"40",
	x"40",
	x"40",
	x"40",

	 -- 385:	0x7F, 0x02, 0x1C, 0x02, 0x7F, 
	x"7F",
	x"02",
	x"1C",
	x"02",
	x"7F",

	 -- 390:	0x7F, 0x04, 0x08, 0x10, 0x7F, 
	x"7F",
	x"04",
	x"08",
	x"10",
	x"7F",

	 -- 395:	0x3E, 0x41, 0x41, 0x41, 0x3E, 
	x"3E",
	x"41",
	x"41",
	x"41",
	x"3E",

	 -- 400:	0x7F, 0x09, 0x09, 0x09, 0x06, 
	x"7F",
	x"09",
	x"09",
	x"09",
	x"06",

	 -- 405:	0x3E, 0x41, 0x51, 0x21, 0x5E, 
	x"3E",
	x"41",
	x"51",
	x"21",
	x"5E",

	 -- 410:	0x7F, 0x09, 0x19, 0x29, 0x46, 
	x"7F",
	x"09",
	x"19",
	x"29",
	x"46",

	 -- 415:	0x26, 0x49, 0x49, 0x49, 0x32, 
	x"26",
	x"49",
	x"49",
	x"49",
	x"32",

	 -- 420:	0x03, 0x01, 0x7F, 0x01, 0x03, 
	x"03",
	x"01",
	x"7F",
	x"01",
	x"03",

	 -- 425:	0x3F, 0x40, 0x40, 0x40, 0x3F, 
	x"3F",
	x"40",
	x"40",
	x"40",
	x"3F",

	 -- 430:	0x1F, 0x20, 0x40, 0x20, 0x1F, 
	x"1F",
	x"20",
	x"40",
	x"20",
	x"1F",

	 -- 435:	0x3F, 0x40, 0x38, 0x40, 0x3F, 
	x"3F",
	x"40",
	x"38",
	x"40",
	x"3F",

	 -- 440:	0x63, 0x14, 0x08, 0x14, 0x63, 
	x"63",
	x"14",
	x"08",
	x"14",
	x"63",

	 -- 445:	0x03, 0x04, 0x78, 0x04, 0x03, 
	x"03",
	x"04",
	x"78",
	x"04",
	x"03",

	 -- 450:	0x61, 0x59, 0x49, 0x4D, 0x43, 
	x"61",
	x"59",
	x"49",
	x"4D",
	x"43",

	 -- 455:	0x00, 0x7F, 0x41, 0x41, 0x41, 
	x"00",
	x"7F",
	x"41",
	x"41",
	x"41",

	 -- 460:	0x02, 0x04, 0x08, 0x10, 0x20, 
	x"02",
	x"04",
	x"08",
	x"10",
	x"20",

	 -- 465:	0x00, 0x41, 0x41, 0x41, 0x7F, 
	x"00",
	x"41",
	x"41",
	x"41",
	x"7F",

	 -- 470:	0x04, 0x02, 0x01, 0x02, 0x04, 
	x"04",
	x"02",
	x"01",
	x"02",
	x"04",

	 -- 475:	0x40, 0x40, 0x40, 0x40, 0x40, 
	x"40",
	x"40",
	x"40",
	x"40",
	x"40",

	 -- 480:	0x00, 0x03, 0x07, 0x08, 0x00, 
	x"00",
	x"03",
	x"07",
	x"08",
	x"00",

	 -- 485:	0x20, 0x54, 0x54, 0x78, 0x40, 
	x"20",
	x"54",
	x"54",
	x"78",
	x"40",

	 -- 490:	0x7F, 0x28, 0x44, 0x44, 0x38, 
	x"7F",
	x"28",
	x"44",
	x"44",
	x"38",

	 -- 495:	0x38, 0x44, 0x44, 0x44, 0x28, 
	x"38",
	x"44",
	x"44",
	x"44",
	x"28",

	 -- 500:	0x38, 0x44, 0x44, 0x28, 0x7F, 
	x"38",
	x"44",
	x"44",
	x"28",
	x"7F",

	 -- 505:	0x38, 0x54, 0x54, 0x54, 0x18, 
	x"38",
	x"54",
	x"54",
	x"54",
	x"18",

	 -- 510:	0x00, 0x08, 0x7E, 0x09, 0x02, 
	x"00",
	x"08",
	x"7E",
	x"09",
	x"02",

	 -- 515:	0x18, 0xA4, 0xA4, 0x9C, 0x78, 
	x"18",
	x"A4",
	x"A4",
	x"9C",
	x"78",

	 -- 520:	0x7F, 0x08, 0x04, 0x04, 0x78, 
	x"7F",
	x"08",
	x"04",
	x"04",
	x"78",

	 -- 525:	0x00, 0x44, 0x7D, 0x40, 0x00, 
	x"00",
	x"44",
	x"7D",
	x"40",
	x"00",

	 -- 530:	0x20, 0x40, 0x40, 0x3D, 0x00, 
	x"20",
	x"40",
	x"40",
	x"3D",
	x"00",

	 -- 535:	0x7F, 0x10, 0x28, 0x44, 0x00, 
	x"7F",
	x"10",
	x"28",
	x"44",
	x"00",

	 -- 540:	0x00, 0x41, 0x7F, 0x40, 0x00, 
	x"00",
	x"41",
	x"7F",
	x"40",
	x"00",

	 -- 545:	0x7C, 0x04, 0x78, 0x04, 0x78, 
	x"7C",
	x"04",
	x"78",
	x"04",
	x"78",

	 -- 550:	0x7C, 0x08, 0x04, 0x04, 0x78, 
	x"7C",
	x"08",
	x"04",
	x"04",
	x"78",

	 -- 555:	0x38, 0x44, 0x44, 0x44, 0x38, 
	x"38",
	x"44",
	x"44",
	x"44",
	x"38",

	 -- 560:	0xFC, 0x18, 0x24, 0x24, 0x18, 
	x"FC",
	x"18",
	x"24",
	x"24",
	x"18",

	 -- 565:	0x18, 0x24, 0x24, 0x18, 0xFC, 
	x"18",
	x"24",
	x"24",
	x"18",
	x"FC",

	 -- 570:	0x7C, 0x08, 0x04, 0x04, 0x08, 
	x"7C",
	x"08",
	x"04",
	x"04",
	x"08",

	 -- 575:	0x48, 0x54, 0x54, 0x54, 0x24, 
	x"48",
	x"54",
	x"54",
	x"54",
	x"24",

	 -- 580:	0x04, 0x04, 0x3F, 0x44, 0x24, 
	x"04",
	x"04",
	x"3F",
	x"44",
	x"24",

	 -- 585:	0x3C, 0x40, 0x40, 0x20, 0x7C, 
	x"3C",
	x"40",
	x"40",
	x"20",
	x"7C",

	 -- 590:	0x1C, 0x20, 0x40, 0x20, 0x1C, 
	x"1C",
	x"20",
	x"40",
	x"20",
	x"1C",

	 -- 595:	0x3C, 0x40, 0x30, 0x40, 0x3C, 
	x"3C",
	x"40",
	x"30",
	x"40",
	x"3C",

	 -- 600:	0x44, 0x28, 0x10, 0x28, 0x44, 
	x"44",
	x"28",
	x"10",
	x"28",
	x"44",

	 -- 605:	0x4C, 0x90, 0x90, 0x90, 0x7C, 
	x"4C",
	x"90",
	x"90",
	x"90",
	x"7C",

	 -- 610:	0x44, 0x64, 0x54, 0x4C, 0x44, 
	x"44",
	x"64",
	x"54",
	x"4C",
	x"44",

	 -- 615:	0x00, 0x08, 0x36, 0x41, 0x00, 
	x"00",
	x"08",
	x"36",
	x"41",
	x"00",

	 -- 620:	0x00, 0x00, 0x77, 0x00, 0x00, 
	x"00",
	x"00",
	x"77",
	x"00",
	x"00",

	 -- 625:	0x00, 0x41, 0x36, 0x08, 0x00, 
	x"00",
	x"41",
	x"36",
	x"08",
	x"00",

	 -- 630:	0x02, 0x01, 0x02, 0x04, 0x02, 
	x"02",
	x"01",
	x"02",
	x"04",
	x"02",

	 -- 635:	0x3C, 0x26, 0x23, 0x26, 0x3C, 
	x"3C",
	x"26",
	x"23",
	x"26",
	x"3C",

	 -- 640:	0x1E, 0xA1, 0xA1, 0x61, 0x12, 
	x"1E",
	x"A1",
	x"A1",
	x"61",
	x"12",

	 -- 645:	0x3A, 0x40, 0x40, 0x20, 0x7A, 
	x"3A",
	x"40",
	x"40",
	x"20",
	x"7A",

	 -- 650:	0x38, 0x54, 0x54, 0x55, 0x59, 
	x"38",
	x"54",
	x"54",
	x"55",
	x"59",

	 -- 655:	0x21, 0x55, 0x55, 0x79, 0x41, 
	x"21",
	x"55",
	x"55",
	x"79",
	x"41",

	 -- 660:	0x22, 0x54, 0x54, 0x78, 0x42, // a-umlaut
	x"22",
	x"54",
	x"54",
	x"78",
	x"42",

	 -- 665:	0x21, 0x55, 0x54, 0x78, 0x40, 
	x"21",
	x"55",
	x"54",
	x"78",
	x"40",

	 -- 670:	0x20, 0x54, 0x55, 0x79, 0x40, 
	x"20",
	x"54",
	x"55",
	x"79",
	x"40",

	 -- 675:	0x0C, 0x1E, 0x52, 0x72, 0x12, 
	x"0C",
	x"1E",
	x"52",
	x"72",
	x"12",

	 -- 680:	0x39, 0x55, 0x55, 0x55, 0x59, 
	x"39",
	x"55",
	x"55",
	x"55",
	x"59",

	 -- 685:	0x39, 0x54, 0x54, 0x54, 0x59, 
	x"39",
	x"54",
	x"54",
	x"54",
	x"59",

	 -- 690:	0x39, 0x55, 0x54, 0x54, 0x58, 
	x"39",
	x"55",
	x"54",
	x"54",
	x"58",

	 -- 695:	0x00, 0x00, 0x45, 0x7C, 0x41, 
	x"00",
	x"00",
	x"45",
	x"7C",
	x"41",

	 -- 700:	0x00, 0x02, 0x45, 0x7D, 0x42, 
	x"00",
	x"02",
	x"45",
	x"7D",
	x"42",

	 -- 705:	0x00, 0x01, 0x45, 0x7C, 0x40, 
	x"00",
	x"01",
	x"45",
	x"7C",
	x"40",

	 -- 710:	0x7D, 0x12, 0x11, 0x12, 0x7D, // A-umlaut
	x"7D",
	x"12",
	x"11",
	x"12",
	x"7D",

	 -- 715:	0xF0, 0x28, 0x25, 0x28, 0xF0, 
	x"F0",
	x"28",
	x"25",
	x"28",
	x"F0",

	 -- 720:	0x7C, 0x54, 0x55, 0x45, 0x00, 
	x"7C",
	x"54",
	x"55",
	x"45",
	x"00",

	 -- 725:	0x20, 0x54, 0x54, 0x7C, 0x54, 
	x"20",
	x"54",
	x"54",
	x"7C",
	x"54",

	 -- 730:	0x7C, 0x0A, 0x09, 0x7F, 0x49, 
	x"7C",
	x"0A",
	x"09",
	x"7F",
	x"49",

	 -- 735:	0x32, 0x49, 0x49, 0x49, 0x32, 
	x"32",
	x"49",
	x"49",
	x"49",
	x"32",

	 -- 740:	0x3A, 0x44, 0x44, 0x44, 0x3A, // o-umlaut
	x"3A",
	x"44",
	x"44",
	x"44",
	x"3A",

	 -- 745:	0x32, 0x4A, 0x48, 0x48, 0x30, 
	x"32",
	x"4A",
	x"48",
	x"48",
	x"30",

	 -- 750:	0x3A, 0x41, 0x41, 0x21, 0x7A, 
	x"3A",
	x"41",
	x"41",
	x"21",
	x"7A",

	 -- 755:	0x3A, 0x42, 0x40, 0x20, 0x78, 
	x"3A",
	x"42",
	x"40",
	x"20",
	x"78",

	 -- 760:	0x00, 0x9D, 0xA0, 0xA0, 0x7D, 
	x"00",
	x"9D",
	x"A0",
	x"A0",
	x"7D",

	 -- 765:	0x3D, 0x42, 0x42, 0x42, 0x3D, // O-umlaut
	x"3D",
	x"42",
	x"42",
	x"42",
	x"3D",

	 -- 770:	0x3D, 0x40, 0x40, 0x40, 0x3D, 
	x"3D",
	x"40",
	x"40",
	x"40",
	x"3D",

	 -- 775:	0x3C, 0x24, 0xFF, 0x24, 0x24, 
	x"3C",
	x"24",
	x"FF",
	x"24",
	x"24",

	 -- 780:	0x48, 0x7E, 0x49, 0x43, 0x66, 
	x"48",
	x"7E",
	x"49",
	x"43",
	x"66",

	 -- 785:	0x2B, 0x2F, 0xFC, 0x2F, 0x2B, 
	x"2B",
	x"2F",
	x"FC",
	x"2F",
	x"2B",

	 -- 790:	0xFF, 0x09, 0x29, 0xF6, 0x20, 
	x"FF",
	x"09",
	x"29",
	x"F6",
	x"20",

	 -- 795:	0xC0, 0x88, 0x7E, 0x09, 0x03, 
	x"C0",
	x"88",
	x"7E",
	x"09",
	x"03",

	 -- 800:	0x20, 0x54, 0x54, 0x79, 0x41, 
	x"20",
	x"54",
	x"54",
	x"79",
	x"41",

	 -- 805:	0x00, 0x00, 0x44, 0x7D, 0x41, 
	x"00",
	x"00",
	x"44",
	x"7D",
	x"41",

	 -- 810:	0x30, 0x48, 0x48, 0x4A, 0x32, 
	x"30",
	x"48",
	x"48",
	x"4A",
	x"32",

	 -- 815:	0x38, 0x40, 0x40, 0x22, 0x7A, 
	x"38",
	x"40",
	x"40",
	x"22",
	x"7A",

	 -- 820:	0x00, 0x7A, 0x0A, 0x0A, 0x72, 
	x"00",
	x"7A",
	x"0A",
	x"0A",
	x"72",

	 -- 825:	0x7D, 0x0D, 0x19, 0x31, 0x7D, 
	x"7D",
	x"0D",
	x"19",
	x"31",
	x"7D",

	 -- 830:	0x26, 0x29, 0x29, 0x2F, 0x28, 
	x"26",
	x"29",
	x"29",
	x"2F",
	x"28",

	 -- 835:	0x26, 0x29, 0x29, 0x29, 0x26, 
	x"26",
	x"29",
	x"29",
	x"29",
	x"26",

	 -- 840:	0x30, 0x48, 0x4D, 0x40, 0x20, 
	x"30",
	x"48",
	x"4D",
	x"40",
	x"20",

	 -- 845:	0x38, 0x08, 0x08, 0x08, 0x08, 
	x"38",
	x"08",
	x"08",
	x"08",
	x"08",

	 -- 850:	0x08, 0x08, 0x08, 0x08, 0x38, 
	x"08",
	x"08",
	x"08",
	x"08",
	x"38",

	 -- 855:	0x2F, 0x10, 0xC8, 0xAC, 0xBA, 
	x"2F",
	x"10",
	x"C8",
	x"AC",
	x"BA",

	 -- 860:	0x2F, 0x10, 0x28, 0x34, 0xFA, 
	x"2F",
	x"10",
	x"28",
	x"34",
	x"FA",

	 -- 865:	0x00, 0x00, 0x7B, 0x00, 0x00, 
	x"00",
	x"00",
	x"7B",
	x"00",
	x"00",

	 -- 870:	0x08, 0x14, 0x2A, 0x14, 0x22, 
	x"08",
	x"14",
	x"2A",
	x"14",
	x"22",

	 -- 875:	0x22, 0x14, 0x2A, 0x14, 0x08, 
	x"22",
	x"14",
	x"2A",
	x"14",
	x"08",

	 -- 880:	0xAA, 0x00, 0x55, 0x00, 0xAA, 
	x"AA",
	x"00",
	x"55",
	x"00",
	x"AA",

	 -- 885:	0xAA, 0x55, 0xAA, 0x55, 0xAA, 
	x"AA",
	x"55",
	x"AA",
	x"55",
	x"AA",

	 -- 890:	0x00, 0x00, 0x00, 0xFF, 0x00, 
	x"00",
	x"00",
	x"00",
	x"FF",
	x"00",

	 -- 895:	0x10, 0x10, 0x10, 0xFF, 0x00, 
	x"10",
	x"10",
	x"10",
	x"FF",
	x"00",

	 -- 900:	0x14, 0x14, 0x14, 0xFF, 0x00, 
	x"14",
	x"14",
	x"14",
	x"FF",
	x"00",

	 -- 905:	0x10, 0x10, 0xFF, 0x00, 0xFF, 
	x"10",
	x"10",
	x"FF",
	x"00",
	x"FF",

	 -- 910:	0x10, 0x10, 0xF0, 0x10, 0xF0, 
	x"10",
	x"10",
	x"F0",
	x"10",
	x"F0",

	 -- 915:	0x14, 0x14, 0x14, 0xFC, 0x00, 
	x"14",
	x"14",
	x"14",
	x"FC",
	x"00",

	 -- 920:	0x14, 0x14, 0xF7, 0x00, 0xFF, 
	x"14",
	x"14",
	x"F7",
	x"00",
	x"FF",

	 -- 925:	0x00, 0x00, 0xFF, 0x00, 0xFF, 
	x"00",
	x"00",
	x"FF",
	x"00",
	x"FF",

	 -- 930:	0x14, 0x14, 0xF4, 0x04, 0xFC, 
	x"14",
	x"14",
	x"F4",
	x"04",
	x"FC",

	 -- 935:	0x14, 0x14, 0x17, 0x10, 0x1F, 
	x"14",
	x"14",
	x"17",
	x"10",
	x"1F",

	 -- 940:	0x10, 0x10, 0x1F, 0x10, 0x1F, 
	x"10",
	x"10",
	x"1F",
	x"10",
	x"1F",

	 -- 945:	0x14, 0x14, 0x14, 0x1F, 0x00, 
	x"14",
	x"14",
	x"14",
	x"1F",
	x"00",

	 -- 950:	0x10, 0x10, 0x10, 0xF0, 0x00, 
	x"10",
	x"10",
	x"10",
	x"F0",
	x"00",

	 -- 955:	0x00, 0x00, 0x00, 0x1F, 0x10, 
	x"00",
	x"00",
	x"00",
	x"1F",
	x"10",

	 -- 960:	0x10, 0x10, 0x10, 0x1F, 0x10, 
	x"10",
	x"10",
	x"10",
	x"1F",
	x"10",

	 -- 965:	0x10, 0x10, 0x10, 0xF0, 0x10, 
	x"10",
	x"10",
	x"10",
	x"F0",
	x"10",

	 -- 970:	0x00, 0x00, 0x00, 0xFF, 0x10, 
	x"00",
	x"00",
	x"00",
	x"FF",
	x"10",

	 -- 975:	0x10, 0x10, 0x10, 0x10, 0x10, 
	x"10",
	x"10",
	x"10",
	x"10",
	x"10",

	 -- 980:	0x10, 0x10, 0x10, 0xFF, 0x10, 
	x"10",
	x"10",
	x"10",
	x"FF",
	x"10",

	 -- 985:	0x00, 0x00, 0x00, 0xFF, 0x14, 
	x"00",
	x"00",
	x"00",
	x"FF",
	x"14",

	 -- 990:	0x00, 0x00, 0xFF, 0x00, 0xFF, 
	x"00",
	x"00",
	x"FF",
	x"00",
	x"FF",

	 -- 995:	0x00, 0x00, 0x1F, 0x10, 0x17, 
	x"00",
	x"00",
	x"1F",
	x"10",
	x"17",

	 -- 1000:	0x00, 0x00, 0xFC, 0x04, 0xF4, 
	x"00",
	x"00",
	x"FC",
	x"04",
	x"F4",

	 -- 1005:	0x14, 0x14, 0x17, 0x10, 0x17, 
	x"14",
	x"14",
	x"17",
	x"10",
	x"17",

	 -- 1010:	0x14, 0x14, 0xF4, 0x04, 0xF4, 
	x"14",
	x"14",
	x"F4",
	x"04",
	x"F4",

	 -- 1015:	0x00, 0x00, 0xFF, 0x00, 0xF7, 
	x"00",
	x"00",
	x"FF",
	x"00",
	x"F7",

	 -- 1020:	0x14, 0x14, 0x14, 0x14, 0x14, 
	x"14",
	x"14",
	x"14",
	x"14",
	x"14",

	 -- 1025:	0x14, 0x14, 0xF7, 0x00, 0xF7, 
	x"14",
	x"14",
	x"F7",
	x"00",
	x"F7",

	 -- 1030:	0x14, 0x14, 0x14, 0x17, 0x14, 
	x"14",
	x"14",
	x"14",
	x"17",
	x"14",

	 -- 1035:	0x10, 0x10, 0x1F, 0x10, 0x1F, 
	x"10",
	x"10",
	x"1F",
	x"10",
	x"1F",

	 -- 1040:	0x14, 0x14, 0x14, 0xF4, 0x14, 
	x"14",
	x"14",
	x"14",
	x"F4",
	x"14",

	 -- 1045:	0x10, 0x10, 0xF0, 0x10, 0xF0, 
	x"10",
	x"10",
	x"F0",
	x"10",
	x"F0",

	 -- 1050:	0x00, 0x00, 0x1F, 0x10, 0x1F, 
	x"00",
	x"00",
	x"1F",
	x"10",
	x"1F",

	 -- 1055:	0x00, 0x00, 0x00, 0x1F, 0x14, 
	x"00",
	x"00",
	x"00",
	x"1F",
	x"14",

	 -- 1060:	0x00, 0x00, 0x00, 0xFC, 0x14, 
	x"00",
	x"00",
	x"00",
	x"FC",
	x"14",

	 -- 1065:	0x00, 0x00, 0xF0, 0x10, 0xF0, 
	x"00",
	x"00",
	x"F0",
	x"10",
	x"F0",

	 -- 1070:	0x10, 0x10, 0xFF, 0x10, 0xFF, 
	x"10",
	x"10",
	x"FF",
	x"10",
	x"FF",

	 -- 1075:	0x14, 0x14, 0x14, 0xFF, 0x14, 
	x"14",
	x"14",
	x"14",
	x"FF",
	x"14",

	 -- 1080:	0x10, 0x10, 0x10, 0x1F, 0x00, 
	x"10",
	x"10",
	x"10",
	x"1F",
	x"00",

	 -- 1085:	0x00, 0x00, 0x00, 0xF0, 0x10, 
	x"00",
	x"00",
	x"00",
	x"F0",
	x"10",

	 -- 1090:	0xFF, 0xFF, 0xFF, 0xFF, 0xFF, 
	x"FF",
	x"FF",
	x"FF",
	x"FF",
	x"FF",

	 -- 1095:	0xF0, 0xF0, 0xF0, 0xF0, 0xF0, 
	x"F0",
	x"F0",
	x"F0",
	x"F0",
	x"F0",

	 -- 1100:	0xFF, 0xFF, 0xFF, 0x00, 0x00, 
	x"FF",
	x"FF",
	x"FF",
	x"00",
	x"00",

	 -- 1105:	0x00, 0x00, 0x00, 0xFF, 0xFF, 
	x"00",
	x"00",
	x"00",
	x"FF",
	x"FF",

	 -- 1110:	0x0F, 0x0F, 0x0F, 0x0F, 0x0F, 
	x"0F",
	x"0F",
	x"0F",
	x"0F",
	x"0F",

	 -- 1115:	0x38, 0x44, 0x44, 0x38, 0x44, 
	x"38",
	x"44",
	x"44",
	x"38",
	x"44",

	 -- 1120:	0xFC, 0x4A, 0x4A, 0x4A, 0x34, // sharp-s or beta
	x"FC",
	x"4A",
	x"4A",
	x"4A",
	x"34",

	 -- 1125:	0x7E, 0x02, 0x02, 0x06, 0x06, 
	x"7E",
	x"02",
	x"02",
	x"06",
	x"06",

	 -- 1130:	0x02, 0x7E, 0x02, 0x7E, 0x02, 
	x"02",
	x"7E",
	x"02",
	x"7E",
	x"02",

	 -- 1135:	0x63, 0x55, 0x49, 0x41, 0x63, 
	x"63",
	x"55",
	x"49",
	x"41",
	x"63",

	 -- 1140:	0x38, 0x44, 0x44, 0x3C, 0x04, 
	x"38",
	x"44",
	x"44",
	x"3C",
	x"04",

	 -- 1145:	0x40, 0x7E, 0x20, 0x1E, 0x20, 
	x"40",
	x"7E",
	x"20",
	x"1E",
	x"20",

	 -- 1150:	0x06, 0x02, 0x7E, 0x02, 0x02, 
	x"06",
	x"02",
	x"7E",
	x"02",
	x"02",

	 -- 1155:	0x99, 0xA5, 0xE7, 0xA5, 0x99, 
	x"99",
	x"A5",
	x"E7",
	x"A5",
	x"99",

	 -- 1160:	0x1C, 0x2A, 0x49, 0x2A, 0x1C, 
	x"1C",
	x"2A",
	x"49",
	x"2A",
	x"1C",

	 -- 1165:	0x4C, 0x72, 0x01, 0x72, 0x4C, 
	x"4C",
	x"72",
	x"01",
	x"72",
	x"4C",

	 -- 1170:	0x30, 0x4A, 0x4D, 0x4D, 0x30, 
	x"30",
	x"4A",
	x"4D",
	x"4D",
	x"30",

	 -- 1175:	0x30, 0x48, 0x78, 0x48, 0x30, 
	x"30",
	x"48",
	x"78",
	x"48",
	x"30",

	 -- 1180:	0xBC, 0x62, 0x5A, 0x46, 0x3D, 
	x"BC",
	x"62",
	x"5A",
	x"46",
	x"3D",

	 -- 1185:	0x3E, 0x49, 0x49, 0x49, 0x00, 
	x"3E",
	x"49",
	x"49",
	x"49",
	x"00",

	 -- 1190:	0x7E, 0x01, 0x01, 0x01, 0x7E, 
	x"7E",
	x"01",
	x"01",
	x"01",
	x"7E",

	 -- 1195:	0x2A, 0x2A, 0x2A, 0x2A, 0x2A, 
	x"2A",
	x"2A",
	x"2A",
	x"2A",
	x"2A",

	 -- 1200:	0x44, 0x44, 0x5F, 0x44, 0x44, 
	x"44",
	x"44",
	x"5F",
	x"44",
	x"44",

	 -- 1205:	0x40, 0x51, 0x4A, 0x44, 0x40, 
	x"40",
	x"51",
	x"4A",
	x"44",
	x"40",

	 -- 1210:	0x40, 0x44, 0x4A, 0x51, 0x40, 
	x"40",
	x"44",
	x"4A",
	x"51",
	x"40",

	 -- 1215:	0x00, 0x00, 0xFF, 0x01, 0x03, 
	x"00",
	x"00",
	x"FF",
	x"01",
	x"03",

	 -- 1220:	0xE0, 0x80, 0xFF, 0x00, 0x00, 
	x"E0",
	x"80",
	x"FF",
	x"00",
	x"00",

	 -- 1225:	0x08, 0x08, 0x6B, 0x6B, 0x08,
	x"08",
	x"08",
	x"6B",
	x"6B",
	x"08",

	 -- 1230:	0x36, 0x12, 0x36, 0x24, 0x36,
	x"36",
	x"12",
	x"36",
	x"24",
	x"36",

	 -- 1235:	0x06, 0x0F, 0x09, 0x0F, 0x06,
	x"06",
	x"0F",
	x"09",
	x"0F",
	x"06",

	 -- 1240:	0x00, 0x00, 0x18, 0x18, 0x00,
	x"00",
	x"00",
	x"18",
	x"18",
	x"00",

	 -- 1245:	0x00, 0x00, 0x10, 0x10, 0x00,
	x"00",
	x"00",
	x"10",
	x"10",
	x"00",

	 -- 1250:	0x30, 0x40, 0xFF, 0x01, 0x01,
	x"30",
	x"40",
	x"FF",
	x"01",
	x"01",

	 -- 1255:	0x00, 0x1F, 0x01, 0x01, 0x1E,
	x"00",
	x"1F",
	x"01",
	x"01",
	x"1E",

	 -- 1260:	0x00, 0x19, 0x1D, 0x17, 0x12,
	x"00",
	x"19",
	x"1D",
	x"17",
	x"12",

	 -- 1265:	0x00, 0x3C, 0x3C, 0x3C, 0x3C,
	x"00",
	x"3C",
	x"3C",
	x"3C",
	x"3C",

	 -- 1270:	0x00, 0x00, 0x00, 0x00, 0x00
	x"00",
	x"00",
	x"00",
	x"00",
	x"00"
);

begin

-- XXX to long par
p0 : process (i_clk,i_reset) is
begin
	if (i_reset = '1') then
		o_character <= (others => '0');
	elsif (rising_edge(i_clk)) then
		o_character <= GLCDFONTC(to_integer(unsigned(i_index)));
	end if;
end  process p0;

--o_character <= GLCDFONTC(to_integer(unsigned(i_index)));

end architecture behavioral_glcdfont;
