--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package p_package is
	constant BYTE_SIZE : integer := 8;
	constant C_CLOCK_COUNTER : integer := 2**16;
end p_package;

package body p_package is
end p_package;
