--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package p_memory_content is

	constant G_BOARD_CLOCK : integer := 50_000_000;
	constant G_BUS_CLOCK : integer := 100_000;
	constant G_ClockDivider : integer := 1000;
	constant G_MemoryAddress : integer := 24;
	constant G_MemoryData : integer := 16;
	subtype MemoryAddress is std_logic_vector(G_MemoryAddress-1 downto 0);
	subtype MemoryDataByte is std_logic_vector(G_MemoryData-1 downto 0);
	constant G_HalfHex : integer := 4;
	constant G_FullHex : integer := G_HalfHex*2;
	constant ROWS : integer := 128;
	constant ROWS_BITS : integer := 7;
	constant COLS_PIXEL : integer := 32;
	constant COLS_PIXEL_BITS : integer := 5;
	constant COLS_BLOCK : integer := 4;
	constant COLS_BLOCK_BITS : integer := 2;
	constant BYTE_BITS : integer := 8;
	constant WORD_BITS : integer := COLS_BLOCK*BYTE_BITS;

	subtype WORD is std_logic_vector(WORD_BITS-1 downto 0);
	type MEMORY is array(ROWS-1 downto 0) of WORD;

	constant memory_content : MEMORY :=
	( -- f              0f              0
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101"),
		("10101010101010101111111111111111"),
		("11111111111111110101010101010101")
		
	);

end p_memory_content;

package body p_memory_content is
end p_memory_content;
