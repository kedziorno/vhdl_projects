library IEEE;
use IEEE.STD_LOGIC_1164.all;
use WORK.p_globals.ALL;

package p_lcd_display is

	type LCDHex is array(G_LCDAnode-1 downto 0) of std_logic_vector(G_HalfHex-1 downto 0);

end p_lcd_display;

package body p_lcd_display is
end p_lcd_display;

