entity n2_core_pll_m1_cust is
port (
vdd_reg : in bit
);
end entity n2_core_pll_m1_cust;
architecture arch of n2_core_pll_m1_cust is
--vss = '1';
begin

end architecture arch;

