entity n2_core_pll_inv_100x_cust is
port (
vdd_reg : in bit;
o : out bit;
i : in bit
);
end entity n2_core_pll_inv_100x_cust;
architecture arch of n2_core_pll_inv_100x_cust is
begin
--wire vss = '0';
o <= not i;
end architecture arch;

